module DT    (input 		     	    clk,
                input			          reset,
                output	            done,
                output			        sti_rd,
                output	    [9:0]	  sti_addr,
                input		    [15:0]	sti_di,
                output	reg		      res_wr,
                output			        res_rd,
                output	reg [13:0]	res_addr,
                output	reg [7:0]	  res_do,
                input		    [7:0]	  res_di   );

  /*----------PARAMETERS--------*/
  parameter  IDLE                = 4'd0;
  parameter  FETCH_ROM_FORWARD   = 4'd1;
  parameter  FETCH_REG_FORWARD   = 4'd2;
  parameter  FORWARD             = 4'd3;
  parameter  BACKWARD_PREPROCESS = 4'd4;
  parameter  FETCH_ROM_BACKWARD  = 4'd5;
  parameter  FETCH_REG_BACKWARD  = 4'd6;
  parameter  BACKWARD            = 4'd7;
  parameter  DONE                = 4'd8;

  //Registers
  reg       eq_reg;
  reg[2:0]  fetch_ram_counter_reg;
  reg[3:0]  current_state,next_state;
  reg[3:0]  counter_reg;
  reg[7:0]  for_back_reg;
  reg[9:0]  rom_addr_index_reg;
  reg[13:0] ram_addr_index_reg;
  reg[15:0] sti_di_reg;

  //flag
  wire  f_r_f_done,forward_done,f_r_f_start;
  wire  f_r_b_done,backward_done,f_r_b_start;
  reg   pad_max_flag;
  wire  skip_f_flag,skip_b_flag,not_object,gt_flag ;

  //wire
  reg  [7:0] min_temp_wire;

  //state
  //wire IDLE_state                 = current_state == IDLE;
  wire FETCH_ROM_FORWARD_state    ;
  wire FETCH_REG_FORWARD_state    ;
  wire FORWARD_state              ;
  wire BACKWARD_PREPROCESS_state  ;
  wire FETCH_ROM_BACKWARD_state   ;
  wire FETCH_REG_BACKWARD_state   ;
  wire BACKWARD_state             ;
  wire DONE_state                 ;

  assign FETCH_ROM_FORWARD_state    = current_state == FETCH_ROM_FORWARD;
  assign FETCH_REG_FORWARD_state    = current_state == FETCH_REG_FORWARD;
  assign FORWARD_state              = current_state == FORWARD;
  assign BACKWARD_PREPROCESS_state  = current_state == BACKWARD_PREPROCESS;
  assign FETCH_ROM_BACKWARD_state   = current_state == FETCH_ROM_BACKWARD;
  assign FETCH_REG_BACKWARD_state   = current_state == FETCH_REG_BACKWARD;
  assign BACKWARD_state             = current_state == BACKWARD;
  assign DONE_state                 = current_state == DONE;

  assign  skip_f_flag = rom_addr_index_reg == 'd0;
  assign  skip_b_flag = rom_addr_index_reg == 'd1023;
  assign  not_object = sti_di_reg[counter_reg] == 0 ;
  assign  gt_flag = for_back_reg >= res_di;

  assign f_r_f_done = (fetch_ram_counter_reg == 'd3 & FETCH_REG_FORWARD_state);
  assign forward_done = (ram_addr_index_reg == 'd16383);
  assign f_r_f_start = (counter_reg == 'd0);

  assign f_r_b_done = (fetch_ram_counter_reg == 'd4 & FETCH_REG_BACKWARD_state);
  assign backward_done = (ram_addr_index_reg == 'd0);
  assign f_r_b_start = (counter_reg == 'd15);

  //sti_addr
  assign sti_addr = sti_rd ? rom_addr_index_reg : 'd0;

  //OUTPUT
  assign done = DONE_state;
  assign sti_rd = FETCH_ROM_FORWARD_state | FETCH_ROM_BACKWARD_state;
  assign res_rd = not_object ? 0 : (FETCH_REG_FORWARD_state | FETCH_REG_BACKWARD_state) ? 1 : 0;

  //res_wr
  always @(negedge clk or negedge reset)
  begin
    if(!reset)
    begin
      res_wr <= 0;
    end
    else
    begin
      res_wr <= FORWARD_state | BACKWARD_state;
    end
  end

  //pad_max_flag
  always @(*)
  begin
    if(ram_addr_index_reg[6:0] == 'd127)
    begin
      pad_max_flag = res_addr[6:0] == 'd0;
    end
    else if(ram_addr_index_reg[6:0] == 'd0)
    begin
      pad_max_flag = res_addr[6:0] == 'd127;
    end
    else if(ram_addr_index_reg[13:7] == 'd127)
    begin
      pad_max_flag = res_addr[13:7] == 'd0;
    end
    else if(ram_addr_index_reg[13:7] == 'd0)
    begin
      pad_max_flag = res_addr[13:7] == 'd127;
    end
    else
    begin
      pad_max_flag = 0;
    end
  end

  //res_addr
  always @(*)
  begin
    if (FETCH_REG_FORWARD_state)
    begin
      case (fetch_ram_counter_reg)
        'd0:
          res_addr = ram_addr_index_reg - 'd129;
        'd1:
          res_addr = ram_addr_index_reg - 'd128;
        'd2:
          res_addr = ram_addr_index_reg - 'd127;
        'd3:
          res_addr = ram_addr_index_reg - 'd1;
        default:
          res_addr = 'd0;
      endcase
    end
    else if(FETCH_REG_BACKWARD_state)
    begin
      case (fetch_ram_counter_reg)
        'd0:
          res_addr = ram_addr_index_reg + 'd1;
        'd1:
          res_addr = ram_addr_index_reg + 'd127;
        'd2:
          res_addr = ram_addr_index_reg + 'd128;
        'd3:
          res_addr = ram_addr_index_reg + 'd129;
        'd4:
          res_addr = ram_addr_index_reg;
        default:
          res_addr = 'd0;
      endcase
    end
    else if(BACKWARD_state | FORWARD_state)
    begin
      res_addr = ram_addr_index_reg;
    end
    else
    begin
      res_addr = 'd0;
    end
  end

  //res_do
  always @(*)
  begin
    if (FORWARD_state)
    begin
      res_do = skip_f_flag ? sti_di_reg[0] : not_object ? 'd0 : for_back_reg + 'd1;
    end
    else if(BACKWARD_state)
    begin
      res_do = skip_b_flag ? sti_di_reg[15] : not_object ? 'd0 : eq_reg ? for_back_reg : for_back_reg + 'd1;
    end
    else
    begin
      res_do = 'd0;
    end
  end

  /*------------CTR---------------*/
  always @(posedge clk or negedge reset)
  begin
    current_state <= !reset ? IDLE : next_state;
  end
  //next_state
  always @(*)
  begin
    case (current_state)
      IDLE:
      begin
        next_state = FETCH_ROM_FORWARD;
      end
      FETCH_ROM_FORWARD:
      begin
        next_state = skip_f_flag ? FORWARD : FETCH_REG_FORWARD;
      end
      FETCH_REG_FORWARD:
      begin
        next_state = not_object ? FORWARD : f_r_f_done ? FORWARD : FETCH_REG_FORWARD;
      end
      FORWARD:
      begin
        next_state = forward_done ? BACKWARD_PREPROCESS : f_r_f_start ? FETCH_ROM_FORWARD : FETCH_REG_FORWARD;
      end
      BACKWARD_PREPROCESS:
      begin
        next_state = FETCH_ROM_BACKWARD;
      end
      FETCH_ROM_BACKWARD:
      begin
        next_state = skip_b_flag ? BACKWARD : FETCH_REG_BACKWARD;
      end
      FETCH_REG_BACKWARD:
      begin
        next_state = not_object ? BACKWARD : f_r_b_done ? BACKWARD : FETCH_REG_BACKWARD;
      end
      BACKWARD:
      begin
        next_state = backward_done ? DONE : f_r_b_start ? FETCH_ROM_BACKWARD : FETCH_REG_BACKWARD ;
      end
      DONE:
      begin
        next_state = IDLE;
      end
      default:
      begin
        next_state = IDLE;
      end
    endcase
  end

  //counter_reg
  always @(posedge clk or negedge reset)
  begin
    if(!reset)
    begin
      counter_reg <= 'd15;
    end
    else if(FORWARD_state)
    begin
      counter_reg <= counter_reg - 'd1;
    end
    else if(BACKWARD_PREPROCESS_state)
    begin
      counter_reg <= 'd0;
    end
    else if(BACKWARD_state)
    begin
      counter_reg <= counter_reg + 'd1;
    end
    else
    begin
      counter_reg <= counter_reg;
    end
  end

  //fetch_ram_counter_reg
  always @(posedge clk or negedge reset)
  begin
    if(!reset)
    begin
      fetch_ram_counter_reg <= 'd0;
    end
    else if(FETCH_REG_FORWARD_state | FETCH_REG_BACKWARD_state)
    begin
      fetch_ram_counter_reg <= fetch_ram_counter_reg + 'd1;
    end
    else if(FORWARD_state | BACKWARD_state)
    begin
      fetch_ram_counter_reg <= 'd0;
    end
    else
    begin
      fetch_ram_counter_reg <= fetch_ram_counter_reg;
    end
  end

  //rom_addr_index_reg
  always @(posedge clk or negedge reset)
  begin
    if(!reset)
    begin
      rom_addr_index_reg <= 'd0;
    end
    else if(FETCH_ROM_FORWARD_state)
    begin
      rom_addr_index_reg <= rom_addr_index_reg + 'd1;
    end
    else if(BACKWARD_PREPROCESS_state)
    begin
      rom_addr_index_reg <= 'd1023;
    end
    else if(FETCH_ROM_BACKWARD_state)
    begin
      rom_addr_index_reg <= rom_addr_index_reg - 'd1;
    end
    else
    begin
      rom_addr_index_reg <= rom_addr_index_reg;
    end
  end

  //ram_addr_index_reg
  always @(posedge clk or negedge reset)
  begin
    if(!reset)
    begin
      ram_addr_index_reg <= 'd0;
    end
    else if(FORWARD_state)
    begin
      ram_addr_index_reg <= ram_addr_index_reg + 'd1;
    end
    else if(BACKWARD_PREPROCESS_state)
    begin
      ram_addr_index_reg <= 'd16383;
    end
    else if(BACKWARD_state)
    begin
      ram_addr_index_reg <= ram_addr_index_reg - 'd1;
    end
    else
    begin
      ram_addr_index_reg <= ram_addr_index_reg;
    end
  end

  //sti_di_reg
  always @(posedge clk or negedge reset)
  begin
    if(!reset)
    begin
      sti_di_reg <= 'd0;
    end
    else if(FETCH_ROM_BACKWARD_state | FETCH_ROM_FORWARD_state)
    begin
      sti_di_reg <= sti_di;
    end
    else
    begin
      sti_di_reg <= sti_di_reg;
    end
  end

  integer i;
  //for_back_reg
  always @(posedge clk or negedge reset)
  begin
    if(!reset)
    begin
      for_back_reg <= 'd0;
    end
    else if(FETCH_REG_FORWARD_state)
    begin
      for_back_reg <= not_object ? 'd0 : min_temp_wire ;
    end
    else if(FETCH_REG_BACKWARD_state)
    begin
      for_back_reg <= not_object ? 'd0 : min_temp_wire ;
    end
    else if(FORWARD_state | BACKWARD_state)
    begin
      for_back_reg <= 'd0;
    end
    else
    begin
      for_back_reg <= for_back_reg;
    end
  end

  //min_temp_wire
  always @(*)
  begin
    if(FETCH_REG_FORWARD_state)
    begin
      case (fetch_ram_counter_reg)
        'd0:
          min_temp_wire = pad_max_flag ? 'd127 : res_di;
        'd1:
          min_temp_wire = pad_max_flag ? for_back_reg : gt_flag ? res_di : for_back_reg;
        'd2:
          min_temp_wire = pad_max_flag ? for_back_reg : gt_flag ? res_di : for_back_reg;
        'd3:
          min_temp_wire = pad_max_flag ? for_back_reg : gt_flag ? res_di : for_back_reg;
        default:
          min_temp_wire = 'd0;
      endcase
    end
    else if(FETCH_REG_BACKWARD_state)
    begin
      case (fetch_ram_counter_reg)
        'd0:
          min_temp_wire = pad_max_flag ? 'd127 : res_di;
        'd1:
          min_temp_wire = pad_max_flag ? for_back_reg : gt_flag ? res_di : for_back_reg;
        'd2:
          min_temp_wire = pad_max_flag ? for_back_reg : gt_flag ? res_di : for_back_reg;
        'd3:
          min_temp_wire = pad_max_flag ? for_back_reg : gt_flag ? res_di : for_back_reg;
        'd4:
          min_temp_wire = gt_flag ? res_di : for_back_reg;
        default:
          min_temp_wire = 'd0;
      endcase
    end
    else
    begin
      min_temp_wire = 'd0;
    end
  end

  //eq_reg
  always @(posedge clk or negedge reset)
  begin
    if(!reset)
    begin
      eq_reg <= 0;
    end
    else if(f_r_b_done)
    begin
      eq_reg <= gt_flag ? 1 : 0;
    end
    else
    begin
      eq_reg <= 0;
    end
  end

endmodule
